package constants is

  constant buswidth : integer := 8;
  constant adr_buswidth : integer := 16;

end constants;
