library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

-- 8x8 16x16 blocks of 8 bit RGB

entity tilemem is

  port(
    clk : in std_logic;
    row_base : in std_logic_vector(2 downto 0);
    row_offset : in std_logic_vector(3 downto 0);
    col_base : in std_logic_vector(2 downto 0);
    col_offset : in std_logic_vector(3 downto 0);
    data_out : out std_logic_vector(7 downto 0));
  
end tilemem;
    
architecture tilemem_behv of tilemem is

  type tilemem_t is array (0 to 16383) of std_logic_vector(7 downto 0);
  signal tilemem : tilemem_t :=(
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00000000",
"11111111", "11111111", "11100000", "11100000", "11100000", "11100000", "11100000", "11100000", "11100000", "11100000", "11100000", "11100000", "11100000", "11111111", "11111111", "00000000",
"00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"00100100", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00100100", "00000000",
"11111111", "11111111", "11111111", "11100000", "11100000", "11100000", "00000000", "00000000", "00000000", "11100000", "11100000", "11100000", "11111111", "11111111", "11111111", "00000000",
"00100100", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "10010010", "00100100", "00000000",
"11100000", "11111111", "11111111", "11111111", "11100000", "00000000", "00000000", "00000000", "00000000", "00000000", "11100000", "11111111", "11111111", "11111111", "11100000", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "10010010", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "10010010", "00100100", "00000000",
"11100000", "11100000", "11111111", "11111111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111111", "11111111", "11100000", "11100000", "00000000",
"00100100", "10010010", "11011011", "00000011", "00000011", "00000011", "00000011", "11111100", "11111100", "00000011", "00000011", "00000000", "11011011", "10010010", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "10010010", "00100100", "00000000",
"11100000", "11100000", "11100000", "00000000", "00000000", "00000000", "00011100", "00000000", "00011100", "00000000", "00000000", "00000000", "11100000", "11100000", "11100000", "00000000",
"00100100", "10010010", "11011011", "00000011", "00000011", "00000011", "00000011", "11111100", "11111100", "00000011", "00000011", "00000000", "11011011", "10010010", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "10010010", "00100100", "00000000",
"11100000", "11100000", "00011100", "00011100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011100", "00011100", "00000000", "11100000", "11100000", "00000000",
"00100100", "10010010", "11011011", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "00000000", "11011011", "10010010", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "10010010", "00100100", "00000000",
"11100000", "00000000", "00011100", "00000000", "00011100", "00000000", "00011100", "00011100", "00011100", "00000000", "00011100", "00000000", "00011100", "00000000", "11100000", "00000000",
"00100100", "10010010", "11011011", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "00000000", "11011011", "10010010", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "10010010", "00100100", "00000000",
"11100000", "00000000", "00011100", "00000000", "00011100", "00000000", "00011100", "00000000", "00011100", "00000000", "00011100", "00000000", "00011100", "00000000", "11100000", "00000000",
"00100100", "10010010", "11011011", "00000011", "00000011", "00000011", "00000011", "11111100", "11111100", "00000011", "00000011", "00000000", "11011011", "10010010", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "10010010", "00100100", "00000000",
"11100000", "00000000", "00011100", "00000000", "00011100", "00000000", "00011100", "00000000", "00011100", "00000000", "00011100", "00000000", "00011100", "00000000", "11100000", "00000000",
"00100100", "10010010", "11011011", "00000011", "00000011", "00000011", "00000011", "11111100", "11111100", "00000011", "00000011", "00000000", "11011011", "10010010", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "10010010", "00100100", "00000000",
"11100000", "11100000", "00011100", "00011100", "00000000", "00000000", "00011100", "00011100", "00011100", "00000000", "00011100", "00011100", "00000000", "11100000", "11100000", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "00000000", "11011011", "10010010", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "10010010", "00100100", "00000000",
"11100000", "11100000", "11100000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11100000", "11100000", "11100000", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "00000000", "11011011", "10010010", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "10010010", "00100100", "00000000",
"11100000", "11100000", "11111111", "11111111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111111", "11111111", "11100000", "11100000", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "00000000", "11011011", "10010010", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "10010010", "00100100", "00000000",
"11100000", "11111111", "11111111", "11111111", "11100000", "00000000", "00000000", "00000000", "00000000", "00000000", "11100000", "11111111", "11111111", "11111111", "11100000", "00000000",
"00100100", "10010010", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "11011011", "10010010", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"10010010", "10010010", "10010010", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "11111111", "11111111", "10010010", "10010010", "10010010", "00000000",
"00100100", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00100100", "00000000",
"11111111", "11111111", "11111111", "11100000", "11100000", "11100000", "00000000", "00000000", "00000000", "11100000", "11100000", "11100000", "11111111", "11111111", "11111111", "00000000",
"00100100", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "00000000",
"00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00000000",
"11111111", "11111111", "11100000", "11100000", "11100000", "11100000", "11100000", "11100000", "11100000", "11100000", "11100000", "11100000", "11100000", "11111111", "11111111", "00000000",
"00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00100100", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00011111", "00011111", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "11111100", "11111100",
"11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100",
"11111100", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100",
"11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100",
"11111100", "11111100", "11111100", "11111100", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "11111100", "11111100", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "11111100", "11111100", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "11111100", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "11111100", "11111100", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "11111100", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "11111100", "11111100", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "11111100", "11111100", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "11111100", "11111100", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100",
"11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100",
"11111100", "11111100", "11111100", "11111100", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "11111100", "11111100",
"11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100", "11111100",
"11111100", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "11111100", "00000000", "11111100", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "11111100", "00000000", "11111100", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "11100011", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000",
"00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000", "00000000"
);
  signal row : std_logic_vector(6 downto 0);
  signal col : std_logic_vector(6 downto 0);
begin

  row <= row_base & row_offset;
  col <= col_base & col_offset;

  process(clk)
  begin
    if rising_edge(clk) then
      data_out <= tilemem(conv_integer(row) * 128 + conv_integer(col));           
    end if;
  end process;
  
end tilemem_behv;
