library ieee;
use work.constants.all;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity micromem is
  port(
		mpc_in : in std_logic_vector(7 downto 0);
		mm_out : out std_logic_vector(1 to 40);
		clk : in std_logic
		);  
end micromem;

architecture micromem_behv of micromem is
  type micromem_type is array (0 to 255) of std_logic_vector(1 to 40);
  signal micromem : micromem_type := ( 																			
-- h�mtfas 0 klar
"1000000000100000010000000000000000000000",
"0000000000100000000000000000000000000000",
"0110100000100000000000000000000000000000",
"0000001100100000000000000000000000000000",
"0000000001000000100000000000000000000000",
-- abs 5 klar
"1000000000100000010000000000000000000000",
"0000000000100000000000000000000000000000",
"0110100000100000100000000000000000000000",
"1000000000100000010000000000000000000000",
"0000000000100000000000000000000000000000",
"0110100000100000000000000000000000000001",
"1000001000100000100000000000000000000000",
"0000000000100000000000000000000000000000",
"0000000010000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- indirekt 15 klar
"1000000000100000010000000000000000000100",  --ar -> hr
"0000000000100000000000000000000000000000",
"0110100000100000100000000000000000000000",
"1000000000100000010000000000000000000000",
"0000000000100000000000000000000000000000",
"0110100000100000000000000000000000000001",
"0000001000100000000000001000000000000000",  --dr -> tr
"0000000000100000000000000010000110000000",  --tr -> ar
"1000001000100000000000000000000000000000",
"0000000000100000000000000011000010000000",  --ar++
"0110100000100000000000000000000000000000",
"1000000000100000000000000000000000001000",
"0000000000100000000000000000000000000000",
"0110100000100000000000000000000000000001",
"1000001010000000100000000000000000000010",  --hr -> ar
-- indexering 30 klar
"0000000000100000000100001000000000000100",
"1000000000100000010000000010000110000000",
"0000000000100000000000000000000000000000",
"0110100000100000100000000000000000000000",
"1000000000100000010000000000000000000000",
"0000000000100000000000000000000000000000",
"0110100000100000000000000000000000000001",
"0000001000100000000000001000000000000000",
"0000000000100000000000000010010010000000",
"1000000000100000000000000000000000001000",
"0000000010000000100000000000000000000010",
-- sj�lvrelativ 41 klar
"1000000000100000010000000000000000000000",
"0000000000100000000000000000000000000000",
"0110100000100000100000000000000000000000",
"1000000000100000010000000000000000000000",
"0000000000100000000000000000000000000000",
"0110100000100000000000000000000000000001",
"0000001000100000000000001000000000000100",
"0000000000100000000000000010000110000000",
"0000000000100000010000001000000000000000",
"0000000000100000000000000010010010000000",
"0000000000100000000000001000000000001000",
"0000000010000000100000000000000000000010",
-- omedelbar 53 klar
"1000000000100000010000000000000000000000",
"0000000010000000100000000000000000000000",
-- underf�rst�dd 55 klar
"0000000010000000000000000000000000000000",
-- LDA 56
"0110100000100000000000000000000000000000",
"0000001000100000000000001000000000000000",
"0000000000100000000000000010000110000000",
"0000000000010000000000000000000001000000",
-- STA 60
"0000010000100000000000000000000000001000",
"0101100000010000000000000000000000000000",
-- ADDA 62                                  
"0110100000100000000000000000000000000000",
"0000001000100000000000001000000000000000",
"0000000000100000000000000010010010000000",
"0000000000010000000000000000000001000000",
-- SUBA 66
"0110100000100000000000000000000000000000",
"0000001000100000000000001000000000000000",
"0000000000100000000000000010001010000000",
"0000000000010000000000000000000001000000",
-- INCA 70
"0000000000100000000000000001000010000000",
"0000000000010000000000000000000001000000",
-- DECA 72
"0000000000100000000000000000100010000000",
"0000000000010000000000000000000001000000",
-- LDX 74                              
"0110100000100000000000000000000000000000",
"0000001000010000001000000000000000000000",
-- STX 76                                
"0000010000100000000100000000000000000000",
"0101100000010000000000000000000000000000",
-- INX 78                        
"0000000000100000000100001000000000000100",
"0000000000100000000000000010000110000000",
"0000000000100000000000000001000010000000",
"0000000000100000001000000000000001001000",
"0000000000010000000000000000000000000010",
-- DEX 83                               
"0000000000100000000100001000000000000100",
"0000000000100000000000000010000110000000",
"0000000000100000000000000000100010000000",
"0000000000100000001000000000000001001000",
"0000000000010000000000000000000000000010",
-- LDS 88                                  HH                             
"0110100000100000000000000000000000000000",
"0000001000010000000010000000000000000000",
-- STS 90
"0000010000100000000000010000000000000000",
"0101100000010000000000000000000000000000",
-- INS 92
"0000000000010000000001000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- DES 97                             
"0000000000010000000000100000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- PUSH 103                   
"1000000000100000000000010000000000000000",  --sp->adr
"0000010000100000000000000000000000001000",  --ar->dr
"0101100000010000000000100000000000000000",  --skriv (sp--)
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- PULL 111                      
"0000000000100000000001000000000000000000",  -- sp++
"1000000000100000000000010000000000000000",  -- sp->adr 
"0110100000100000000000000000000000000000",  -- l�s
"0000001000100000000000001000000000000000",  -- dr->tr
"0000000000100000000000000010000110000000",  -- tr->ar
"0000000000010000000000000000000001000000",  -- ar->sr (mpc = 0)
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- JMP 122
"0000000000011000000000000100000000000000",                              
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- JPMN 127                                    
"0000000000010110000000000100000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- JMPZ 133
"0000000000010101000000000100000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- JSR 139                                   
"1000000000100000000000010000000000000000",
"0000010000100000010000000000000000000000",
"0101100000011000000000100100000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- RTS 146
"1000000000100000000000010000000000000000",
"0110100000100000000000000000000000000000",
"0000001000011000000001000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- HH 153 klar
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- LSR 155 klar
"0000000000100000000000000001000110000000",
"0000000000010000000000000000000001000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- LSL 160 klar
"0000000000100000000000000001001010000000",
"0000000000010000000000000000000001000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- ASR 165 klar
"0000000000100000000000000001010010000000",
"0000000000010000000000000000000001000000",
"0000000000100000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- ASL 170 klar
"0000000000000000000000000001100010000000",
"0000000000010000000000000000000001000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- AND 175
"0110100000100000000000000000000000000000",
"0000001000100000000000001000000000000000",
"0000000000100000000000000011110010000000",
"0000000000010000000000000000000000000000",
"0000000000000000000000000000000000000000",
-- CMP 180
"0000000000100000000000000000000000000000",
"0110100000100000000000000000000000000100",
"0000001000100000000000001000000000000000",
"0000000000100000000000000010001010000000",
"0000000000010000000000000000000001000010",
-- LDA16 185
"0110100000100000000000000000000000000000",
"1000000000100000010000000000000000000000",
"0000000000100000000000000000000000000000",
"0110100000100000100000000000000000000001",
"0000001000100000000000001000000000000000",
"0000000000100000000000000010000110000000",
"0000000000010000000000000000000001000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000",
--STA16 195 (endast absolut)
"0000000000100000000000000000000000000100", --ar->hr
"0000001000100000000000001001000110000000",  --LSRx8 (dr->tr)
"0000000000100000000000000001000110000000",
"0000000000100000000000000001000110000000",
"0000000000100000000000000001000110000000",
"0000000000100000000000000001000110000000",
"0000000000100000000000000001000110000000",
"0000000000100000000000000001000110000000",
"0000000000100000000000000001000110000000",
"0000010000100000000000000010000110001000",  --ar->dr, tr->ar
"0101100000100000000000000001000010000000",  --skriv
"1000000000100000000000000000000000001000",  --ar->adr
"0000000000100000000000000000000000000010",  --hr->ar
"0000010000100000000000000000000000001000",  --ar->dr
"0101100000010000000000000000000000000000",  --skriv
--ADDA16 210
"0000000000100000000000000000000000000000",
"0110100000100000000000000000000000000000",  --l�s (pc++)
"1000000000100000010000000000000000000000",  --pc->adr
"0000000000100000000000000000000000000000",  --v�nta
"0110100000100000100000000000000000000001",  --l�s (skifta)
"0000001000100000000000001000000000000000",  --dr->tr
"0000000000100000000000000010010010000000",  --add
"0000000000100000000000000000000000000000",
"0000000000010000000000000000000001000000",  --ar->sr

others => "0000000000000000000000000000000000000000");

begin
	       mm_out <= micromem(conv_integer(mpc_in));
end micromem_behv;
