package constants is

  constant bus_width : integer := 8;

end constants;
