package constants is

  constant buswidth : integer := 8;

end constants;
