package constants is

  constant buswidth : integer := 16;
  constant adr_buswidth : integer := 16;

end constants;
