library IEEE;
use work.constants.all;
use IEEE.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity primmem is    
   port (
	 clk : in std_logic;
     adr_bus : in std_logic_vector(15 downto 0);
	 data_bus_in : in std_logic_vector(7 downto 0);
	 data_bus_out : out std_logic_vector(7 downto 0);
	 read_signal : in std_logic;
	 write_signal : in std_logic);
end primmem;

architecture primmem_behv of primmem is

type primmem_type is array (0 to 4095) of std_logic_vector(7 downto 0);
  signal primmem : primmem_type := (
-- S�tt stackpekare. 0
    
"01010100",-- 0:                             -- LDS omedelbar
"00001111",-- 1:
"11111111",-- 2:                 -- #4095


-- Initialisera variabler.

-- Bomber minus flaggor 3
"00000100",-- 3:                             -- LDA omedelbar
"00101000",-- 4:                             -- #40
"00001000",-- 5:                             -- STA absolut
"00001100",                             -- 6:
"00011011",-- 7:                 -- $3099

-- Global end game flagga 8
"00000100",-- 8:                             -- LDA omedelbar
"00000000",-- 9:                             -- #0
"00001000",-- 10:                             -- STA absolut
"00001100",                             -- 11:
"00011010",-- 12:                 -- $3098

-- Initialisera spelplan. 28
    
"00000100",-- 13:                             -- LDA omedelbar
"01000000",-- 14:                             -- #64
"00110100",-- 15:                             -- LDX omedelbar
"11111111",-- 16:                             -- #255
"00001010",-- 17:                             -- STA indexerad
"00001100",                             -- 18:
"00011100",-- 19:                 -- #3100
"01001101",-- 20:                             -- DEX
"10001011",-- 21:                             -- JMPN relativ
"00000000",                             -- 22:
"00000100",-- 23:                 -- #4
"10000011",-- 24:                             -- JMP relativ
"11111111",                             -- 25:
"11110111",-- 26:                 -- #-9

    
-- Placera minor. 42

"00110100",-- 27:                             -- LDX omedelbar
"00101000",-- 28:                             -- #40
-- H�mta slumptal.
"00000000",-- 29:                             -- LDA abs
"00100000",                             -- 30:
"00000001",-- 31:                 -- $8193
-- Skapa x-offset. 47
"11010100",-- 32:                             -- AND omedelbar
"00001111",-- 33:                             -- #15
"00001000",-- 34:                             -- STA absolut
-- Spara x-offset i 3000. 
"00001011",                             -- 35:
"10111000",-- 36:                 -- $3000
-- Skapa y-offset. 52
"00000000",-- 37:                             -- LDA abs
"00100000",                             -- 38:
"00000001",-- 39:                 -- $8193
"11010100",-- 40:                             -- AND omedelbar
"00001111",-- 41:                             -- #15
"10111101",-- 42:                             -- LSL
"10111101",-- 43:                             -- LSL
"10111101",-- 44:                             -- LSL
"10111101",-- 45:                             -- LSL
-- L�gg ihop x och y-offset. 61
"00010000",-- 46:                             -- ADD absolut
"00001011",                             -- 47:
"10111000",-- 48:                 -- $3000
-- L�gg till konstant (pekare in i spelplansdatastrukturen).
"11110100",-- 49:                             -- ADD16 omedelbar
"00001100",                             -- 50:
"00011100",-- 51:                 -- #3100
-- Spara adress i 3001.
"11101000",-- 52:                             -- STA16 absolut
"00001011",                             -- 53:
"10111001",-- 54:                 -- $3001
-- Ladda A med v�rdet f�r en osynlig mina.
"00000100",-- 55:                             -- LDA omedelbar
"01001011",-- 56:                             -- #11
-- Kolla om en mina redan ligger p� den platsen.
"11011001",-- 57:                             -- CMP indirekt
"00001011",                             -- 58:
"10111001",-- 59:                 -- $3001
-- B�rja om isf. 75
"10010011",-- 60:                             -- JMPZ relativ
"11111111",                             -- 61:
"11011111",-- 62:                 -- #-33
-- Spara minan i datastrukturen.
"00001001",-- 63:                             -- STA indirekt
"00001011",                             -- 64:
"10111001",-- 65:                 -- $3001
-- R�kna ner och b�rja om. 81
"01001101",-- 66:                             -- DEX
"10010011",-- 67:                             -- JMPZ
"00000000",                             -- 68:
"00000101",-- 69:                 -- #5
"10000011",-- 70:                             -- JMP -43
"11111111",                             -- 71:
"11010101",                             -- 72:
"10101101",-- 73:                             -- HH


-- Generera siffror. 89

"00110100",-- 74:                             -- LDX omedelbar
"11111111",-- 75:                             -- #255
-- Kolla mina och slut.
"00000010",-- 76:                             -- LDA indexerad
"00001100",                             -- 77:
"00011100",-- 78:                 -- #3100
"11010100",-- 79:                             -- AND omedelbar
"00001111",-- 80:                             -- #15
"11011100",-- 81:                             -- CMP omedelbar
"00001011",-- 82:                             -- #11
"10010011",-- 83:                             -- JMPZ
"00000000",                             -- 84:
"00001000",                             -- 85:
"01001101",-- 86:                             -- DEX
"10001011",-- 87:                             -- JMPN SLUT
"00000000",                             -- 88:
"01110100",                             -- 89:
"10000011",-- 90:                             -- JMP b�rjan
"11111111",                             -- 91:
"11110000",                             -- 92:
-- Initiera y- och x-till�gg. 108
"11100100",-- 93:                             -- LDA16
"11111111",                             -- 94:
"11110000",-- 95:                 -- -16
"11101000",-- 96:                             -- STA16
"00001011",                             -- 97:
"10111000",-- 98:                 -- $3000
"11100100",-- 99:                             -- LDA16
"11111111",                             -- 100:
"11111111",-- 101:                 -- -1
"11101000",-- 102:                             -- STA16
"00001011",                             -- 103:
"10111010",-- 104:                 -- $3002
-- y-bounds 120
"00111000",-- 105:                             -- STX
"00001011",                             -- 106:
"10111100",-- 107:                 -- $3004
"00000000",-- 108:                             -- LDA
"00001011",                             -- 109:
"10111100",-- 110:                 -- $3004
"11010100",-- 111:                             -- AND
"11110000",                             -- 112:
"11000000",-- 113:                             -- ADD16ABSOLUT
"00001011",                             -- 114:
"10111000",-- 115:                 -- $3000
"10001011",-- 116:                             -- JMPN
"00000000",                             -- 117:
"01000111",-- 118:                 -- 71 
"10110101",-- 119:                             -- LSR
"11011100",-- 120:                             -- CMP
"10000000",-- 121:                             -- #128
"10010011",-- 122:                             -- JMPZ
"00000000",                             -- 123:
"01000001",-- 124:                 -- 65
"10111101",-- 125:                             -- LSL
"00001000",-- 126:                             -- STA
"00001011",                             -- 127:
"10111101",-- 128:                 -- $3005
-- x-bounds 144
"00000000",-- 129:                             -- LDA
"00001011",                             -- 130:
"10111100",-- 131:                 -- $3004
"11010100",-- 132:                             -- AND
"00001111",-- 133:                             -- #15
"11000000",-- 134:                             -- ADD16ABSOLUT
"00001011",                             -- 135:
"10111010",-- 136:                 -- $3002
"10001011",-- 137:                             -- JMPN
"00000000",                             -- 138:
"00100011",-- 139:                 -- 35
"11011100",-- 140:                             -- CMP
"00010000",-- 141:                             -- #16
"10010011",-- 142:                             -- JMPZ
"00000000",                             -- 143:
"00011110",-- 144:                 -- 30
"00001000",-- 145:                              --STA
"00001011",                             -- 146:
"10111110",-- 147:                 -- $3006
"00010000",-- 148:                             -- ADD
"00001011",                             -- 149:
"10111101",-- 150:                 -- $3005
"11110100",-- 151:                             -- ADD16
"00001100",                             -- 152:
"00011100",-- 153:                 -- #3100
"11101000",-- 154:                             -- STA16ABSOLUT
"00001011",                             -- 155:
"10111111",-- 156:                 -- $3007
"00000001",-- 157:                             -- LDA
"00001011",                             -- 158:
"10111111",-- 159:                 -- $3007
"11010100",-- 160:                             -- AND
"00001111",-- 161:                             -- #15
"11011100",-- 162:                             -- CMP
"00001011",-- 163:                             -- mina
"10010011",-- 164:                             -- JMPZ
"00000000",                             -- 165:
"00001000",-- 166:                 -- 8
"00000001",-- 167:                             -- LDA
"00001011",                             -- 168:
"10111111",-- 169:                 -- $3007
"00100101",-- 170:                             -- INC
"00001001",-- 171:                             -- STA
"00001011",                             -- 172:
"10111111",-- 173:                 -- $3007
--n�sta x 189
"11111000",-- 174:                             -- LDA16ABSOLUT
"00001011",                             -- 175:
"10111010",-- 176:                 -- $3002
"00100101",-- 177:                             -- INC
"11101000",-- 178:                             -- STA16ABSOLUT
"00001011",                             -- 179:
"10111010",-- 180:                 -- $3002
"11011100",-- 181:                             -- CMP
"00000010",-- 182:                             -- #2
"10010011",-- 183:                             -- JMPZ n�sta y
"00000000",                             -- 184:
"00000100",-- 185:                 -- 4
"10000011",-- 186:                             -- JMP x_bound
"11111111",                             -- 187:
"11000101",-- 188:                 -- -59
--n�sta y 204
"11111000",-- 189:                             -- LDA16ABSOLUT
"00001011",                             -- 190:
"10111000",-- 191:                 -- $3000
"00010100",-- 192:                             -- ADD
"00010000",-- 193:                             -- #16
"11101000",-- 194:                             -- STA16ABSOLUT
"00001011",                             -- 195:
"10111000",-- 196:                 -- $3000
"11011100",-- 197:                             -- CMP
"00100000",-- 198:                             -- #32
"10010011",-- 199:                             -- JMPZ 
"11111111",                             -- 200:
"10001101",-- 201:                 -- -115
"10000011",-- 202:                             -- JMP (y-bounds)
"11111111",                             -- 203:
"10010111",-- 204:                 -- -105


-- Main loop. 

"10011011",-- 205:                             -- JSR rita spelplan
"00000000",                             -- 206:
"00001101",-- 207:                 -- #13
"10011011",-- 208:                             -- JSR statusrad
"00000000",                             -- 209:
"01100101",-- 210:                 -- 101
"10011011",-- 211:                             -- JSR mushantering
"00000000",                             -- 212:
"10110010",-- 213:                 -- #178
"10011011",-- 214:                             -- JSR End-Game 
"00000010",                             -- 215:
"01000101",-- 216:                 -- #508+3+51 
"10000011",-- 217:                             -- JMP
"11111111",                             -- 218:
"11110010",-- 219:                 -- #-14


-- Rita spelplan. 235

-- V�nta p� VSYNC.
"00000000",-- 220:                             -- LDA absolut
"00100000",                             -- 221:
"00001001",-- 222:                 -- $8201
"11010100",-- 223:                             -- AND omedelbar
"00000001",-- 224:                             -- #1
"10010011",-- 225:                             -- JMPZ relativ
"11111111",                             -- 226:
"11111001",-- 227:                 -- #-7
-- Ladda indexr�knaren.
"00110100",-- 228:                             -- LDX omedelbar
"11111111",-- 229:                             -- #255
"00111000",-- 230:                             -- STX absolut
"00001011",                             -- 231:
"10111000",-- 232:                 -- $3000
"00000000",-- 233:                             -- LDA absolut
"00001011",                             -- 234:
"10111000",-- 235:                 -- $3000
-- x-offset 251
"11010100",-- 236:                             -- AND omedelbar
"00001111",-- 237:                             -- #15
"00001000",-- 238:                             -- STA absolut
"00001011",                             -- 239:
"10111001",-- 240:                 -- $3001
-- y-offset 256
"00000000",-- 241:                             -- LDA absolut
"00001011",                             -- 242:
"10111000",-- 243:                 -- $3000
"11010100",-- 244:                             -- AND omedelbar
"11110000",-- 245:                             -- #240
"10111101",-- 246:                             -- LSL underf�rst�dd
"10111101",-- 247:                             -- LSL underf�rst�dd
"00010000",-- 248:                             -- ADD absolut
"00001011",                             -- 249:
"10111001",-- 250:                 -- $3001
-- L�gg till konstant till adressen.
"11110100",-- 251:                             -- ADD16 omedelbar
"00010001",           --600                  -- 252:
"11001100",-- 253:                 -- #4096
-- Spara adress till grafikminnet i 3002.
"11101000",-- 254:                             -- STA16 absolut
"00001011",                             -- 255:
"10111010",-- 256:                 -- $3002
-- Kolla om vi ska rita en flagga.
"00000010",-- 257:                             -- LDA indexerad
"00001100",                             -- 258:
"00011100",-- 259:                 -- #3100
"11010100",-- 260:                             -- AND omedelbar
"01000000",-- 261:                             -- #64
"10010011",-- 262:                             -- JMPZ relativ
"00000000",                             -- 263:
"00010110",-- 264:                 -- #22
-- Kolla om vi ska rita ett osynligt block. 281
"00000010",-- 265:                             -- LDA indexerad
"00001100",                             -- 266:
"00011100",-- 267:                 -- #3100
"11010100",-- 268:                             -- AND omedelbar
"10000000",-- 269:                             -- #128
"10010011",-- 270:                             -- JMPZ relativ
"00000000",                             -- 271:
"00011010",-- 272:                 -- #26
-- Rita synligt block. 288
"00000010",-- 273:                             -- LDA indexerad
"00001100",                             -- 274:
"00011100",-- 275:                 -- #3100
"00001001",-- 276:                             -- STA indirekt
"00001011",                             -- 277:
"10111010",-- 278:                 -- $3002
"01001101",-- 279:                             -- DEX underf�rst�dd
"10001011",-- 280:                             -- JMPN relativ
"00000000",                             -- 281:
"00011100",-- 282:                 -- #28
"10000011",-- 283:                             -- JMP relativ
"11111111",                             -- 284:
"11001001",-- 285:                 -- #-55
-- Rita flagga. 301
"00000100",-- 286:                             -- LDA omedelbar
"00001100",-- 287:                             -- #12
"00001001",-- 288:                             -- STA indirekt
"00001011",                             -- 289:
"10111010",-- 290:                 -- $3002
"01001101",-- 291:                             -- DEX underf�rst�dd
"10001011",-- 292:                             -- JMPN relativ
"00000000",                             -- 293:
"00010000",-- 294:                 -- #16
"10000011",-- 295:                             -- JMP relativ
"11111111",                             -- 296:
"10111101",                             -- 297:
-- Rita osynligt block. 313
"00000100",-- 298:                             -- LDA omedelbar
"00001010",-- 299:                             -- #10
"00001001",-- 300:                             -- STA indirekt
"00001011",                             -- 301:
"10111010",-- 302:                 -- $3002
"01001101",-- 303:                             -- DEX underf�rst�dd
"10001011",-- 304:                             -- JMPN relativ
"00000000",                             -- 305:
"00000100",                             -- 306:
"10000011",-- 307:                             -- JMP relativ
"11111111",                             -- 308:
"10110001",                             -- 309:
"10100101",-- 310:                             -- RTS


-- 101 fr�n hopp i mainanrop
-- Rita statusrad. 326

"00000000",-- 311:                             -- LDA
"00100000",                             -- 312:
"00001000",-- 313:                 -- $8200
"00010100",-- 314:                             -- ADD omedelbar
"00010000",-- 315:                             -- #16
"00001000",-- 316:                             -- STA
"00010001",                             -- 317:
"10010001",-- 318:                 -- $4497
"00000000",-- 319:                             -- LDA
"00100000",                             -- 320:
"00000111",-- 321:                 -- $8199
"00010100",-- 322:                             -- ADD omedelbar
"00010000",-- 323:                             -- #16
"00001000",-- 324:                             -- STA
"00010001",                             -- 325:
"10010010",-- 326:                 -- $4498
"00000000",-- 327:                             -- LDA
"00100000",                             -- 328:
"00000110",-- 329:                 -- $8198
"00010100",-- 330:                             -- ADD omedelbar
"00010000",-- 331:                             -- #16
"00001000",-- 332:                             -- STA
"00010001",                             -- 333:
"10010011",-- 334:                 -- $4499
"00000100",-- 335:                             -- LDA
"00001010",-- 336:                             -- #10
"00001000",-- 337:                             -- STA
"00001011",                             -- 338:
"11101010",-- 339:                 -- $3050 -- n�mnare
"00000000",-- 340:                             -- LDA
"00001100",                             -- 341:
"00011011",-- 342:                 -- $3099
"00001000",-- 343:                             -- STA
"00001011",                             -- 344:
"11101011",-- 345:                 -- $3051 -- t�ljare
"10011011",-- 346:                             -- JSR division
"00000001",                             -- 347:
"11111010",-- 348:                 -- #18
"00000000",-- 349:                             -- LDA
"00001011",                             -- 350:
"11101100",-- 351:                 -- $3052 kvot
"00010100",-- 352: 500                             -- ADD omedelbar
"00010000",-- 353:                             -- #16
"00001000",-- 354:                             -- STA
"00010001",                             -- 355:
"10010101",-- 356:                 -- $4501
"00000000",-- 357:                             -- LDA
"00001011",                             -- 358:
"11101101",-- 359:                 -- $3053 rest
"00010100",-- 360:                             -- ADD omedelbar
"00010000",-- 361:                             -- #16
"00001000",-- 362:                             -- STA
"00010001",                             -- 363:
"10010110",-- 364:                 -- $4502
"10100101",-- 365:                             -- RTS


-- 155 fr�n main-funktionen
-- Division 381
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",
"00000110",


-- Mushantering 

-- Spara xpos
"00000000",-- 391:                             -- LDA absolut
"00100000",                             -- 392:
"00000011",-- 393:                 -- $8195
"00001000",-- 394:                             -- STA absolut
"00001011",                             -- 395:
"10111000",-- 396:                 -- $3000
-- Spara ypos 412
"00000000",-- 397:                             -- LDA absolut
"00100000",                             -- 398:
"00000100",-- 399:                 -- $8196
"00001000",-- 400:                             -- STA absolut
"00001011",                             -- 401:
"10111001",-- 402:                 -- $3001
-- R�kna ut adress 418
"01011101",-- 403:                             -- LSLx4
"00010000",-- 404:                             -- ADD absolut
"00001011",                             -- 405:
"10111000",-- 406:                 -- $3000
"11110100",-- 407:                             -- ADD16 omedelbar
"00001100",                             -- 408:
"00011100",-- 409:                 -- #3100
"11101000",-- 410:                             -- STA16 absolut
"00001011",                             -- 411:
"10111011",-- 412:                 -- $3003
-- Hantera klick 428
"00000000",-- 413:                             -- LDA absolut
"00100000",                             -- 414:
"00000010",-- 415:                 -- klick $8194
"00001000",-- 416:                             -- STA absolut
"00001011",                             -- 417:
"10111010",-- 418:                 -- $3002
"11010100",-- 419:                             -- AND omedelbar
"10000000",-- 420:                             -- #128
"10010011",-- 421:                             -- JMPZ hoppa till h�gerklick-hantering
"00000000",                             -- 422:
"00101100",-- 423:                 -- 44
-- Kolla om cellen �r synlig 439
"00000001",-- 424:                             -- LDA indirekt
"00001011",                             -- 425:
"10111011",-- 426:                 -- $3003
"11010100",-- 427:                             -- AND omedelbar
"10000000",-- 428:                             -- #128 
"10010011",-- 429:                             -- JMPZ hoppa �ver rts
"00000000",                             -- 430:
"00000010",-- 431:                 -- #2
"10100101",-- 432:                             -- RTS (g� ur)
-- Kolla om cellen �r flaggad 448
"00000001",-- 433:                             -- LDA indirekt
"00001011",                             -- 434:
"10111011",-- 435:                 -- $3003
"11010100",-- 436:                             -- AND omedelbar
"01000000",-- 437:                             -- #64
"10010011",-- 438:                             -- JMPZ g� ur
"11111111",                             -- 439:
"11111000",-- 440:                 -- #-8
-- Kolla om cellen �r en mina 456
"00000001",-- 441:                             -- LDA indirekt
"00001011",                             -- 442:
"10111011",-- 443:                 -- $3003
"11011100",-- 444:                             -- CMP omedelbar
"01001011",-- 445:                             -- #75 (kolla om mina)
"10010011",-- 446:                             -- JMPZ end-game
"00000000",                             -- 447:
"01110100",-- 448:                 -- #46+51
"00110100",-- 449:                             -- LDX omedelbar
"00000000",-- 450:                             -- #0
-- Cellen �r tom eller numrerad, starta flood-fill 466
"00000000",-- 451:                             -- LDA absolut
"00001011",            --400                 -- 452:
"10111000",-- 453:                 -- $3000 x-pos
"00001010",-- 454:                             -- STA index
"00000111",                             -- 455:
"11010001",-- 456:                 -- $2001
"00000000",-- 457:                             -- LDA absolut
"00001011",                             -- 458:
"10111001",-- 459:                 -- $3001 y-pos
"00001010",-- 460:                             -- STA index
"00000111",                             -- 461:
"11010000",-- 462:                 -- $2000
"10011011",-- 463:                             -- JSR (Flood Fill) 
"00000000",                             -- 464:
"01101001",-- 465:                 -- #32+3+51
"10100101",-- 466:                             -- RTS
-- H�gerklick 482
-- Kolla om h�gerklick
"00000000",-- 467:                             -- LDA absolut
"00001011",                             -- 468:
"10111010",-- 469:                 -- $3002 klick-info
"11010100",-- 470:                             -- AND omedelbar
"00000001",-- 471:                             -- #1 h�gerklick
"10010011",-- 472:                             -- JMPZ hoppa tll rts
"11111111",                             -- 473:
"11111000",-- 474:                 -- #-8
-- NYTT SKIT Kolla om det g�tt en sekund sen sista h�gerklicket
-- Kolla sekund
"00000000",-- 475:                             -- LDA absolut
"00100000",                             -- 476:
"00000110",-- 477:                  -- $8198
"11011000",-- 478:                             -- CMP absolut
"00001100",                             -- 479:
"00001010",-- 480:                  -- $3082
"10010011",-- 481:                             -- JMPZ tiotal
"00000000",                             -- 482:
"00000100",-- 483:                  -- #4
"10000011",-- 484:                             -- JMP forts�tt
"00000000",                             -- 485:
"00010110",-- 486:                  -- #22
-- Kolla tiotals sekunder 13
"00000000",-- 487:                             -- LDA absolut
"00100000",                             -- 488:
"00000111",-- 489:                  -- $8199
"11011000",-- 490:                             -- CMP absolut
"00001100",                             -- 491:
"00001001",-- 492:                  -- $3081
"10010011",-- 493:                             -- JMPZ hundratal
"00000000",                             -- 494:
"00000100",-- 495:                  -- #4
"10000011",-- 496:                             -- JMP forts�tt
"00000000",                             -- 497:
"00001010",-- 498:                  -- #10
-- Kolla hundratals sekunder 25
"00000000",-- 499:                             -- LDA absolut
"00100000",                             -- 500:
"00001000",-- 501:                  -- $8200
"11011000",-- 502:                             -- CMP absolut
"00001100",                             -- 503:
"00001000",-- 504:                  -- $3080
"10010011",-- 505:                             -- JMPZ avsluta
"00000000",                             -- 506:
"00011011",-- 507:                  -- #28
-- Spara ny tid f�r senaste h�gerklick 34
"00000000",-- 508:                             -- LDA absolut
"00100000",                             -- 509:
"00000110",-- 510:                  -- $8198
"00001000",-- 511:                             -- STA absolut
"00001100",                             -- 512:
"00001010",-- 513:                  -- $3082
"00000000",-- 514:                             -- LDA absolut
"00100000",                             -- 515:
"00000111",-- 516:                  -- $8199
"00001000",-- 517:  --301                           -- STA absolut
"00001100",                             -- 518:
"00001001",-- 519:                  -- $3081
"00000000",-- 520:                             -- LDA absolut
"00100000",                             -- 521:
"00001000",-- 522:                  -- $8200
"00001000",-- 523:                             -- STA absolut
"00001100",                             -- 524:
"00001000",-- 525:                  -- $3080
-- SLUT NYTT SKIT 51 l�ng
-- Kolla om cellen �r synlig 490 + 51
"00000001",-- 526:                             -- LDA indirekt
"00001011",                             -- 527:
"10111011",-- 528:                 -- $3003 spelplanscell
"11010100",-- 529:                             -- AND omedelbar
"10000000",-- 530:                             -- #128 en rad borttagen
"10010011",-- 531:                             -- JMPZ hoppa �ver rts
"00000000",                             -- 532:
"00000010",-- 533:                 -- #2
"10100101",-- 534:                             -- RTS
-- Cellen �r osynlig, toggla flagga 500 --
"00000001",-- 535:                             -- LDA indirekt
"00001011",                             -- 536:
"10111011",-- 537:                 -- 3003 spelplanscell (v�rdet f�rst�rt
                                        -- av and) 3 nya rader
"10101100",-- 538:                             -- XOR omedelbar
"01000000",-- 539:                             -- #64 toggla flagga
"00001001",-- 540:                             -- STA indirekt
"00001011",                             -- 541:
"10111011",-- 542:                 -- $3003 spelplanscell
"11010100",-- 543:                             -- AND omedelbar
"01000000",-- 544:                             -- #64
"10010011",-- 545:                             -- JMPZ s�nk flaggr�knaren
"00000000",                             -- 546:
"00001001",-- 547:                 -- #9
"00000000",-- 548:                             -- LDA absolut
"00001100",                             -- 549:
"00011011",-- 550:                 -- $3099
"00100101",-- 551:                             -- INCA
"00001000",-- 552:  300                           -- STA absolut
"00001100",                             -- 553:
"00011011",-- 554:                 -- $3099
"10100101",-- 555:                             -- RTS
"00000000",-- 556:                             -- LDA absolut
"00001100",                             -- 557:
"00011011",-- 558:                 -- $3099
"00101101",-- 559:                             -- DECA
"00001000",-- 560:                             -- STA absolut
"00001100",                             -- 561:
"00011011",-- 562:                 -- $3099
"10100101",-- 563:                             -- RTS
-- End-game, s�tt end-game flagga i minnet
"00000100",-- 564:                             -- LDA omedelbar
"00000001",-- 565:                             -- #1 
"00001000",-- 566:                             -- STA absolut
"00001100",                             -- 567:
"00011010",-- 568:                 -- $3098 game over flagga
"10100101",-- 569:   --53                          -- RTS


-- Flood fill 515
-- H�mta ypos
"00000010",-- 570:                             -- LDA index
"00000111",                             -- 571:
"11010000",-- 572:                 -- $2000
-- Kolla om ypos �r giltig
"11010100",-- 573:                             -- AND omedelbar
"11110000",-- 574:                             -- #240
"10010011",-- 575:                             -- JMPZ
"00000000",                             -- 576:
"00000010",-- 577:                 -- #2
-- Hoppar ur rekursionen 523
"10100101",-- 578:                             -- RTS
-- H�mta xpos
"00000010",-- 579:                             -- LDA index
"00000111",                             -- 580:
"11010001",-- 581:                 -- $2001
-- Kolla om xpos �r giltig
"11010100",-- 582:                             -- AND omedelbar
"11110000",-- 583:                             -- #240
"10010011",-- 584:                             -- JMPZ
"00000000",                             -- 585:
"00000010",-- 586:                 -- #2
-- Hoppa ur rekursionen 532
"10100101",-- 587:                             -- RTS
-- R�kna ut adress
"00000010",-- 588:                             -- LDA8 indexerad
"00000111",                             -- 589:
"11010000",-- 590:                 -- $2000
"01011101",-- 591:                             -- LSLx4
"00010010",-- 592:                             -- ADD index
"00000111",                             -- 593:
"11010001",-- 594:                 -- $2001
"11110100",-- 595:                             -- ADD16 omedelbar
"00001100",                             -- 596:
"00011100",-- 597:                 -- #3100
"11101000",-- 598:                             -- STA16 absolut
"00001011",                             -- 599:
"10111010",-- 600:                 -- $3002
-- H�mta cellen 546
"00000001",-- 601:                             -- LDA indirekt
"00001011",                             -- 602:
"10111010",-- 603:                 -- $3002
-- Kolla om cellen �r flaggad
"11010100",-- 604:                             -- AND
"01000000",-- 605:                             -- #64
-- Hoppa ur om cellen �r flaggad 550
"10010011",-- 606:                             -- JMPZ 
"00000000",                             -- 607:
"00001001",-- 608:                 -- #9
-- H�mta cellen igen
"00000001",-- 609:                             -- LDA indirekt
"00001011",                             -- 610:
"10111010",-- 611:                 -- $3002
-- Kolla om cellen �r synlig
"11010100",-- 612:                             -- AND omedelbar
"10000000",-- 613:                             -- #128
-- Hoppa till 'g�r cellen synlig'
"10010011",-- 614:                             -- JMPZ
"00000000",                             -- 615:
"00000010",-- 616:                 -- #2
-- Hoppa ur rekursionen 562
"10100101",-- 617:     --401                        -- RTS
-- G�r cellen synlig
"00000001",-- 618:                             -- LDA indirekt
"00001011",                             -- 619:
"10111010",-- 620:                 -- $3002
"11001100",-- 621:                             -- OR omedelbar
"10000000",-- 622:                             -- #128
"00001001",-- 623:                             -- STA indirekt
"00001011",                             -- 624:
"10111010",-- 625:                 -- $3002
-- Kolla om cellen �r en nolla 571
"11010100",-- 626:                             -- AND omedelbar
"00001111",-- 627:                             -- #15
-- Hoppa till rekursivt anrop
"10010011",-- 628:                             -- JMPZ
"00000000",                             -- 629:
"00000010",-- 630:                 -- 2
-- Hoppa ur rekursionen
"10100101",-- 631:                             -- RTS
-- Rekursivt anrop
-- Nord 577
-- Spara ny xpos
"00000010",-- 632:                             -- LDA indexerad
"00000111",                             -- 633:
"11010001",-- 634:                 -- $2001
"00001010",-- 635:                             -- STA indexerad
"00000111",                             -- 636:
"11010011",-- 637:                 -- $2003
-- Spara ny ypos
"00000010",-- 638:                             -- LDA indexerad
"00000111",                             -- 639:
"11010000",-- 640:                 -- $2000
"00101101",-- 641:                             -- DECA
"00001010",-- 642:                             -- STA indexerad
"00000111",                             -- 643:
"11010010",-- 644:                 -- $2002
-- �ka indexeringen 590
"01000101",-- 645:                             -- INX
"01000101",-- 646:                             -- INX
-- Starta om algoritm
"10011011",-- 647:                             -- JSR
"11111111",                             -- 648:
"10110001",-- 649:                 -- #-79
"01001101",-- 650:                             -- DEX
"01001101",-- 651:                             -- DEX
-- NYTT SKIT
-- Nordost 597
-- Spara ny xpos
"00000010",-- 652:    200                         -- LDA indexerad
"00000111",                             -- 653:
"11010001",-- 654:                 -- $2001
"00100101",-- 655:                             -- INCA
"00001010",-- 656:                             -- STA indexerad
"00000111",                             -- 657:
"11010011",-- 658:                 -- $2003
-- Spara ny ypos 604
"00000010",-- 659:                              -- LDA indexerad
"00000111",                             -- 660:
"11010000",-- 661:                 -- $2000
"00101101",-- 662:                             -- DECA
"00001010",-- 663:                             -- STA indexerad
"00000111",                             -- 664:
"11010010",-- 665:                 -- $2002
-- �ka indexeringen
"01000101",-- 666:                             -- INX
"01000101",-- 667:                             -- INX
-- Starta om algoritm
"10011011",-- 668:                             -- JSR
"11111111",                             -- 669:
"10011100",-- 670:                 -- #-100
"01001101",-- 671:                             -- DEX
"01001101",-- 672:                             -- DEX
-- Ost 618
-- Spara ny xpos
"00000010",-- 673:                             -- LDA indexerad
"00000111",                             -- 674:
"11010001",-- 675:                 -- $2001
"00100101",-- 676:                             -- INCA
"00001010",-- 677:                             -- STA indexerad
"00000111",                             -- 678:
"11010011",-- 679:                 -- $2003
-- Spara ny ypos
"00000010",-- 680:                             -- LDA indexerad
"00000111",                             -- 681:
"11010000",-- 682:                 -- $2000
"00001010",-- 683:                             -- STA indexerad
"00000111",                             -- 684:
"11010010",-- 685:                 -- $2002
-- �ka indexeringen
"01000101",-- 686:                             -- INX
"01000101",-- 687:                             -- INX
-- Starta om algoritm
"10011011",-- 688:                             -- JSR
"11111111",                             -- 689:
"10001000",-- 690:                 -- #-120
"01001101",-- 691:                             -- DEX
"01001101",-- 692:                             -- DEX
-- Sydost 638
-- Spara ny xpos
"00000010",-- 693:                             -- LDA indexerad
"00000111",                             -- 694:
"11010001",-- 695:                 -- $2001
"00100101",-- 696:                             -- INCA
"00001010",-- 697:                             -- STA indexerad
"00000111",                             -- 698:
"11010011",-- 699:                 -- $2003
-- Spara ny ypos
"00000010",-- 700:                             -- LDA indexerad
"00000111",                             -- 701:
"11010000",-- 702:                 -- $2000
"00100101",-- 703:                             -- INCA
"00001010",-- 704:                             -- STA indexerad
"00000111",                             -- 705:
"11010010",-- 706:                 -- $2002
-- �ka indexeringen
"01000101",-- 707:                             -- INX
"01000101",-- 708:                             -- INX
-- Starta om algoritm
"10011011",-- 709:                             -- JSR
"11111111",                             -- 710:
"01110011",-- 711:                 -- #-141
"01001101",-- 712:                             -- DEX
"01001101",-- 713:--97(98?)                             -- DEX
-- Syd 659
-- Spara ny xpos
"00000010",-- 714:                             -- LDA indexerad
"00000111",                             -- 715:
"11010001",-- 716:                 -- $2001
"00001010",-- 717:                             -- STA indexerad
"00000111",                             -- 718:
"11010011",-- 719:                 -- $2003
-- Spara ny ypos
"00000010",-- 720:                             -- LDA indexerad
"00000111",                             -- 721:
"11010000",-- 722:                 -- $2000
"00100101",-- 723:                             -- INCA
"00001010",-- 724:                             -- STA indexerad
"00000111",                             -- 725:
"11010010",-- 726:                 -- $2002
-- �ka indexeringen
"01000101",-- 727:                             -- INX
"01000101",-- 728:                             -- INX
-- Starta om algoritm 674
"10011011",-- 729:                             -- JSR
"11111111",                             -- 730:
"01011111",-- 731:                 -- #-161
"01001101",-- 732:                             -- DEX
"01001101",-- 733:                             -- DEX
-- Sydv�st 679
-- Spara ny xpos
"00000010",-- 734:                             -- LDA indexerad
"00000111",                             -- 735:
"11010001",-- 736:                 -- $2001
"00101101",-- 737:                             -- DECA
"00001010",-- 738:                             -- STA indexerad
"00000111",                             -- 739:
"11010011",-- 740:                 -- $2003
-- Spara ny ypos
"00000010",-- 741:                             -- LDA indexerad
"00000111",                             -- 742:
"11010000",-- 743:                 -- $2000
"00100101",-- 744:                             -- INCA
"00001010",-- 745:                             -- STA indexerad
"00000111",                             -- 746:
"11010010",-- 747:                 -- $2002
-- �ka indexeringen
"01000101",-- 748:                             -- INX
"01000101",-- 749:                             -- INX
-- Starta om algoritm
"10011011",-- 750:                             -- JSR
"11111111",                             -- 751:
"01001010",-- 752: 100                 -- #-182
"01001101",-- 753:                             -- DEX
"01001101",-- 754:                             -- DEX
-- V�st 700
-- Spara ny xpos
"00000010",-- 755:                             -- LDA indexerad
"00000111",                             -- 756:
"11010001",-- 757:                 -- $2001
"00101101",-- 758:                             -- DECA
"00001010",-- 759:                             -- STA indexerad
"00000111",                             -- 760:
"11010011",-- 761:                 -- $2003
-- Spara ny ypos
"00000010",-- 762:                             -- LDA indexerad
"00000111",                             -- 763:
"11010000",-- 764:                 -- $2000
"00001010",-- 765:                             -- STA indexerad
"00000111",                             -- 766:
"11010010",-- 767:                 -- $2002
-- �ka indexeringen
"01000101",-- 768:                             -- INX
"01000101",-- 769:                             -- INX
-- Starta om algoritm
"10011011",-- 770:                             -- JSR
"11111111",                             -- 771:
"00110110",-- 772:                 -- #-202
"01001101",-- 773:                             -- DEX
"01001101",-- 774:                             -- DEX
-- Nordv�st 720
-- Spara ny xpos
"00000010",-- 775:                             -- LDA indexerad
"00000111",                             -- 776:
"11010001",-- 777:                 -- $2001
"00101101",-- 778:                             -- DECA
"00001010",-- 779:                             -- STA indexerad
"00000111",                             -- 780:
"11010011",-- 781:                 -- $2003
-- Spara ny ypos
"00000010",-- 782:                             -- LDA indexerad
"00000111",                             -- 783:
"11010000",-- 784:                 -- $2000
"00101101",-- 785:                             -- DECA
"00001010",-- 786:                             -- STA indexerad
"00000111",                             -- 787:
"11010010",-- 788:                 -- $2002
-- �ka indexeringen 734
"01000101",-- 789:                             -- INX
"01000101",-- 790:                             -- INX
-- Starta om algoritm
"10011011",-- 791:                             -- JSR
"11111111",                             -- 792:
"00100001",-- 793:                 -- #-223
"01001101",-- 794:                             -- DEX
"01001101",-- 795:                             -- DEX
-- SLUT NYTT SKIT 741
"10100101",-- 796:                             -- RTS


-- End Game 742+51
-- Kolla om spelet �r vunnet
"00110100",                             -- LDX omedelbar
"11111111",                             -- #255
"00000010",                             -- LDA indexerad
"00001100",
"00011100",                             -- #3100
"11010100",                             -- AND omedelbar
"00001011",                             -- #mina
"11011100",                             -- CMP omedelbar
"00001011",                             -- #mina
"10010011",                             -- JMPZ mina
"00000000",
"00001001",                             -- 12
"00000010",                             -- LDA indexerad
"00001100",
"00011100",                             -- #3100
"11010100",                             -- AND omedelbar
"10000000",                             -- #128
"10010011",                             -- JMPZ avsluta 
"00000000",
"00001000",                             -- 8
"01001101",                             -- DEX
"10001011",                             -- JMPN vunnit
"00000000",
"00011110",                             -- 30
"10000011",                             -- JMP
"11111111",
"11101000",                             -- -24
-- Ladda global End-game-flagga
"00000000",-- 797:                         -- LDA absolut
"00001100",                             -- 798:
"00011010",-- 799:                 -- $3098
"11011100",-- 800:                             -- CMP
"00000001",-- 801:                             -- #1
"10010011",-- 802:                             -- JMPZ
"00000000",                             -- 803:
"00000010",-- 804:                 -- #2
"10100101",-- 805:                             -- RTS
"00110100",-- 806:                             -- LDX omedelbar
"11111111",-- 807:                             -- #255
-- H�mta spelcell
"00000010",-- 808:                             -- LDA indexerad
"00001100",                             -- 809:
"00011100",-- 810:                 -- #3100
-- G�r cellen synlig
"11001100",-- 811:                             -- OR omedelbar
"10000000",-- 812:                             -- #128
-- Spara cellen
"00001010",-- 813:                             -- STA indexerad
"00001100",                             -- 814:
"00011100",-- 815:                 -- #3100
-- B�rja om
"01001101",-- 816:                             -- DEX
"10001011",-- 817:                             -- JMPN relativ
"00000000",                             -- 818:
"00000100",-- 819:                 -- #4
"10000011",-- 820:                             -- JMP relativ
"11111111",                             -- 821:
"11110010",-- 822:                 -- #-14
-- Rita ut spelplan
"10011011",-- 823:                             -- JSR 
"11111101",                             -- 824:
"10001000",-- 825:                 -- -607
-- HALT i Tengils namn
"00000111",                             -- 826:


-- Division

"00110100",-- 366:                             -- LDX
"00000000",-- 367:                             -- #0
"00000000",-- 368:                             -- LDA
"00001011",                             -- 369:
"11101011",-- 370:                 -- $3051 -- t�ljare
"00011000",-- 371:                             -- SUB
"00001011",                             -- 372:
"11101010",-- 373:                 -- $3050 -- n�mnare
"10001011",-- 374:                             -- JMPN
"00000000",                             -- 375:
"00000101",-- 376:                 -- 5
"01000101",-- 377:                             -- INX
"10000011",-- 378:                             -- JMP
"11111111",                             -- 379:
"11110111",-- 380:                 -- -9
"00010000",                             -- 381:
                             -- ADD
"00001011",                             -- 382:
"11101010",-- 383:                 -- $3050 -- n�mnare
"00001000",-- 384:                             -- STA
"00001011",                             -- 385:
"11101101",-- 386:                 -- $3053 rest
"00111000",-- 387:                             -- STX
"00001011",                             -- 388:
"11101100",-- 389:                 -- $3052 kvot
"00000000",                             -- LDA absolut
"00001011",
"11101100",                             -- $3052
"11010100",                             -- AND absolut
"11111000",                             -- #248
"10010011",                             -- JMPZ
"00000000",
"00001001",
"00000100",                             -- LDA omedelbar
"00000000",                             -- #0
"00001000",                             -- STA absolut
"00001011",
"11101100",                             -- $3052
"00001000",                             -- STA absolut
"00001011",
"11101101",                             -- $3053
"10100101",-- 390:                             -- RTS

 
others =>"00000000"
);

begin
  process(clk)
    begin
      if rising_edge(clk) then
          data_bus_out <= primmem(conv_integer(adr_bus));
        if write_signal ='1' then
          primmem(conv_integer(adr_bus)) <= data_bus_in;
      end if;
    end if;
    end process;            
end primmem_behv;

