library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

-- 8x8 16x16 blocks of 8 bit RGB

entity micromem is

  port(
		mpc_in : in std_logic_vector(7 downto 0);
		mm_out : out std_logic_vector(1 to 39)
		);
  
end micromem;

architecture micromem_behv of micromem is

  type micromem_type is array (0 to 255) of std_logic_vector(1 to 39);
  signal micromem : micromem_type := ( 																			-- 4x64
"100000000010000001000000000000000000000", "011010000100000000000000000000000000000", "000000110010000000000000000000000000000", "000000000100000010000000000000000000000",	-- hämtfas
"100000000010000001000000000000000000000", "011010000010000000000000000000000000000", "100000101000000100000000000000000000000", -- abs
"100000000010000001000000000000000000000", "011010000010000000000000000000000000000", "100000100010000000000000000000000000000", 
"011010000010000000000000000000000000000", "100000101000000010000000000000000000000", -- indirekt
"000000000010000000010000100000000000000", "100000000000000001000000001000010000000", "011010000010000000000000000000000000000", 
"000000100010000000000000100000000000000", "000000000010000000000000001001001000000", "100000000010000000000000000000000000100", "000000001000000010000000000000000000000", -- indexering
"100000000010000001000000000000000000000", "011010000010000010000000000000000000000", "000000100010000000000000100000000000000", "000000000010000000000000001000011000000", 
"000000000010000001000000100000000000000", "000000000010000000000000001001001000000", "000000000010000000000000100000000000100", "000000001000000000000000000000000000000", -- självrelativ
"100000000010000001000000000000000000000", "000000001000000010000000000000000000000", -- omedelbar
"000000001000000000000000000000000000000", --underförstådd
"011010000010000000000000000000000000000", "000000100010000000000010000000000000000", "000000000010000000000000001000011000000", "000000000001000000000000000000000100000", -- ladda ackumulator
"000001000010000000000000000000000000100", "010110000001000000000000000000000000000", -- STA
"011010000010000000000000000000000000000", "000000100010000000000000100000000000000", "000000000010000000000000001001001000000", "000000000001000000000000000000000100000", -- add ackumulator
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000010000000010000100000000000000", "000000000010000000000000001000011000000", "000000000010000000000000000100001000000", "000000000010000000100000000000000100100",
"000000000001000000000000000000000000000", -- INX 
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"100000000010000000000001000000000000000", "000001000010000000000000000000000000100", "010110000001000000000010000000000000000", -- PUSH
"000000000010000000000100000000000000000", "100000000010000000000001000000000000000", "011010000010000000000000000000000000000", 
"000000100010000000000000100000000000000", "000000000010000000000000001000011000000", "000000000001000000000000000000000100000", -- Pull
"000000000001100000000000010000000000000", -- JMP
"000000000001011000000000010000000000000", -- JMPN
"000000000001010100000000010000000000000", -- JMPZ
"100000000010000000000010000000000000000", "000001000010000001000000000000000000000", "010110000001100000000010010000000000000", -- JSR
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
"000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000", "000000000000000000000000000000000000000",
);
begin
	mm_out <= micromem(mpc_in);
	
end tilemem_behv;
